// pc2_perm.v - DES Permuted Choice 2 (PC-2)
module pc2_perm(
    input  [55:0] cd56,    // {C, D}
    output [47:0] k48
);
    assign k48 = {
        cd56[56-14], cd56[56-17], cd56[56-11], cd56[56-24], cd56[56-1],  cd56[56-5],
        cd56[56-3],  cd56[56-28], cd56[56-15], cd56[56-6],  cd56[56-21], cd56[56-10],
        cd56[56-23], cd56[56-19], cd56[56-12], cd56[56-4],  cd56[56-26], cd56[56-8],
        cd56[56-16], cd56[56-7],  cd56[56-27], cd56[56-20], cd56[56-13], cd56[56-2],
        cd56[56-41], cd56[56-52], cd56[56-31], cd56[56-37], cd56[56-47], cd56[56-55],
        cd56[56-30], cd56[56-40], cd56[56-51], cd56[56-45], cd56[56-33], cd56[56-48],
        cd56[56-44], cd56[56-49], cd56[56-39], cd56[56-56], cd56[56-34], cd56[56-53],
        cd56[56-46], cd56[56-42], cd56[56-50], cd56[56-36], cd56[56-29], cd56[56-32]
    };
endmodule

// ---- S-Boxes (FIPS 46-3) ----
module des_sboxes(input [47:0] in48, output [31:0] out32);
    function [3:0] s1; input [5:0] b; integer r,c; begin
        r = {b[5],b[0]}; c = b[4:1];
        case (r)
          0: case(c)
            0: s1=14; 1: s1=4;  2: s1=13; 3: s1=1;  4: s1=2;  5: s1=15; 6: s1=11; 7: s1=8;
            8: s1=3;  9: s1=10; 10: s1=6; 11: s1=12;12: s1=5; 13: s1=9; 14: s1=0;  15: s1=7;
          endcase
          1: case(c)
            0: s1=0;  1: s1=15; 2: s1=7;  3: s1=4;  4: s1=14; 5: s1=2;  6: s1=13; 7: s1=1;
            8: s1=10; 9: s1=6;  10:s1=12; 11:s1=11;12: s1=9; 13: s1=5; 14: s1=3;  15: s1=8;
          endcase
          2: case(c)
            0: s1=4;  1: s1=1;  2: s1=14; 3: s1=8;  4: s1=13; 5: s1=6;  6: s1=2;  7: s1=11;
            8: s1=15; 9: s1=12; 10:s1=9;  11:s1=7; 12: s1=3; 13: s1=10;14: s1=5;  15: s1=0;
          endcase
          default: case(c)
            0: s1=15; 1: s1=12; 2: s1=8;  3: s1=2;  4: s1=4;  5: s1=9;  6: s1=1;  7: s1=7;
            8: s1=5;  9: s1=11; 10:s1=3;  11:s1=14;12: s1=10;13: s1=0; 14: s1=6;  15: s1=13;
          endcase
        endcase
    end endfunction

    function [3:0] s2; input [5:0] b; integer r,c; begin
        r={b[5],b[0]}; c=b[4:1];
        case(r)
          0: case(c)
            0: s2=15;1: s2=1; 2: s2=8; 3: s2=14;4: s2=6; 5: s2=11;6: s2=3; 7: s2=4;
            8: s2=9; 9: s2=7;10: s2=2; 11: s2=13;12:s2=12;13:s2=0;14:s2=5;15:s2=10;
          endcase
          1: case(c)
            0: s2=3; 1: s2=13;2: s2=4; 3: s2=7; 4: s2=15;5: s2=2; 6: s2=8; 7: s2=14;
            8: s2=12;9: s2=0;10: s2=1; 11: s2=10;12:s2=6; 13:s2=9;14:s2=11;15:s2=5;
          endcase
          2: case(c)
            0: s2=0; 1: s2=14;2: s2=7; 3: s2=11;4: s2=10;5: s2=4; 6: s2=13;7: s2=1;
            8: s2=5; 9: s2=8;10: s2=12;11: s2=6; 12:s2=9; 13:s2=3; 14:s2=2; 15:s2=15;
          endcase
          default: case(c)
            0: s2=13;1: s2=8; 2: s2=10;3: s2=1; 4: s2=3; 5: s2=15;6: s2=4; 7: s2=2;
            8: s2=11;9: s2=6;10: s2=7; 11: s2=12;12:s2=0; 13:s2=5; 14:s2=14;15:s2=9;
          endcase
        endcase
    end endfunction

    function [3:0] s3; input [5:0] b; integer r,c; begin
        r={b[5],b[0]}; c=b[4:1];
        case(r)
          0: case(c)
            0:s3=10;1:s3=0; 2:s3=9; 3:s3=14;4:s3=6; 5:s3=3; 6:s3=15;7:s3=5;
            8:s3=1; 9:s3=13;10:s3=12;11:s3=7; 12:s3=11;13:s3=4;14:s3=2;15:s3=8;
          endcase
          1: case(c)
            0:s3=13;1:s3=7; 2:s3=0; 3:s3=9; 4:s3=3; 5:s3=4; 6:s3=6; 7:s3=10;
            8:s3=2; 9:s3=8;10:s3=5; 11:s3=14;12:s3=12;13:s3=11;14:s3=15;15:s3=1;
          endcase
          2: case(c)
            0:s3=13;1:s3=6; 2:s3=4; 3:s3=9; 4:s3=8; 5:s3=15;6:s3=3; 7:s3=0;
            8:s3=11;9:s3=1;10:s3=2; 11:s3=12;12:s3=5; 13:s3=10;14:s3=14;15:s3=7;
          endcase
          default: case(c)
            0:s3=1; 1:s3=10;2:s3=13;3:s3=0; 4:s3=6; 5:s3=9; 6:s3=8; 7:s3=7;
            8:s3=4; 9:s3=15;10:s3=14;11:s3=3; 12:s3=11;13:s3=5; 14:s3=2; 15:s3=12;
          endcase
        endcase
    end endfunction

    function [3:0] s4; input [5:0] b; integer r,c; begin
        r={b[5],b[0]}; c=b[4:1];
        case(r)
          0: case(c)
            0:s4=7; 1:s4=13;2:s4=14;3:s4=3; 4:s4=0; 5:s4=6; 6:s4=9; 7:s4=10;
            8:s4=1; 9:s4=2; 10:s4=8; 11:s4=5; 12:s4=11;13:s4=12;14:s4=4; 15:s4=15;
          endcase
          1: case(c)
            0:s4=13;1:s4=8; 2:s4=11;3:s4=5; 4:s4=6; 5:s4=15;6:s4=0; 7:s4=3;
            8:s4=4; 9:s4=7; 10:s4=2; 11:s4=12;12:s4=1; 13:s4=10;14:s4=14;15:s4=9;
          endcase
          2: case(c)
            0:s4=10;1:s4=6; 2:s4=9; 3:s4=0; 4:s4=12;5:s4=11;6:s4=7; 7:s4=13;
            8:s4=15;9:s4=1;10:s4=3; 11:s4=14;12:s4=5; 13:s4=2; 14:s4=8; 15:s4=4;
          endcase
          default: case(c)
            0:s4=3; 1:s4=15;2:s4=0; 3:s4=6; 4:s4=10;5:s4=1; 6:s4=13;7:s4=8;
            8:s4=9; 9:s4=4; 10:s4=5; 11:s4=11;12:s4=12;13:s4=7; 14:s4=2; 15:s4=14;
          endcase
        endcase
    end endfunction

    function [3:0] s5; input [5:0] b; integer r,c; begin
        r={b[5],b[0]}; c=b[4:1];
        case(r)
          0: case(c)
            0:s5=2; 1:s5=12;2:s5=4; 3:s5=1; 4:s5=7; 5:s5=10;6:s5=11;7:s5=6;
            8:s5=8; 9:s5=5; 10:s5=3; 11:s5=15;12:s5=13;13:s5=0;14:s5=14;15:s5=9;
          endcase
          1: case(c)
            0:s5=14;1:s5=11;2:s5=2; 3:s5=12;4:s5=4; 5:s5=7; 6:s5=13;7:s5=1;
            8:s5=5; 9:s5=0; 10:s5=15;11:s5=10;12:s5=3; 13:s5=9; 14:s5=8; 15:s5=6;
          endcase
          2: case(c)
            0:s5=4; 1:s5=2; 2:s5=1; 3:s5=11;4:s5=10;5:s5=13;6:s5=7; 7:s5=8;
            8:s5=15;9:s5=9;10:s5=12;11:s5=5; 12:s5=6; 13:s5=3; 14:s5=0; 15:s5=14;
          endcase
          default: case(c)
            0:s5=11;1:s5=8; 2:s5=12;3:s5=7; 4:s5=1; 5:s5=14;6:s5=2; 7:s5=13;
            8:s5=6; 9:s5=15;10:s5=0; 11:s5=9; 12:s5=10;13:s5=4; 14:s5=5; 15:s5=3;
          endcase
        endcase
    end endfunction

    function [3:0] s6; input [5:0] b; integer r,c; begin
        r={b[5],b[0]}; c=b[4:1];
        case(r)
          0: case(c)
            0:s6=12;1:s6=1; 2:s6=10;3:s6=15;4:s6=9; 5:s6=2; 6:s6=6; 7:s6=8;
            8:s6=0; 9:s6=13;10:s6=3; 11:s6=4; 12:s6=14;13:s6=7; 14:s6=5; 15:s6=11;
          endcase
          1: case(c)
            0:s6=10;1:s6=15;2:s6=4; 3:s6=2; 4:s6=7; 5:s6=12;6:s6=9; 7:s6=5;
            8:s6=6; 9:s6=1; 10:s6=13;11:s6=14;12:s6=0; 13:s6=11;14:s6=3; 15:s6=8;
          endcase
          2: case(c)
            0:s6=9; 1:s6=14;2:s6=15;3:s6=5; 4:s6=2; 5:s6=8; 6:s6=12;7:s6=3;
            8:s6=7; 9:s6=0; 10:s6=4; 11:s6=10;12:s6=1; 13:s6=13;14:s6=11;15:s6=6;
          endcase
          default: case(c)
            0:s6=4; 1:s6=3; 2:s6=2; 3:s6=12;4:s6=9; 5:s6=5; 6:s6=15;7:s6=10;
            8:s6=11;9:s6=14;10:s6=1; 11:s6=7; 12:s6=6; 13:s6=0; 14:s6=8; 15:s6=13;
          endcase
        endcase
    end endfunction

    function [3:0] s7; input [5:0] b; integer r,c; begin
        r={b[5],b[0]}; c=b[4:1];
        case(r)
          0: case(c)
            0:s7=4; 1:s7=11;2:s7=2; 3:s7=14;4:s7=15;5:s7=0; 6:s7=8; 7:s7=13;
            8:s7=3; 9:s7=12;10:s7=9; 11:s7=7; 12:s7=5; 13:s7=10;14:s7=6; 15:s7=1;
          endcase
          1: case(c)
            0:s7=13;1:s7=0; 2:s7=11;3:s7=7; 4:s7=4; 5:s7=9; 6:s7=1; 7:s7=10;
            8:s7=14;9:s7=3;10:s7=5; 11:s7=12;12:s7=2; 13:s7=15;14:s7=8; 15:s7=6;
          endcase
          2: case(c)
            0:s7=1; 1:s7=4; 2:s7=11;3:s7=13;4:s7=12;5:s7=3; 6:s7=7; 7:s7=14;
            8:s7=10;9:s7=15;10:s7=6; 11:s7=8; 12:s7=0; 13:s7=5; 14:s7=9; 15:s7=2;
          endcase
          default: case(c)
            0:s7=6; 1:s7=11;2:s7=13;3:s7=8; 4:s7=1; 5:s7=4; 6:s7=10;7:s7=7;
            8:s7=9; 9:s7=5; 10:s7=0; 11:s7=15;12:s7=14;13:s7=2; 14:s7=3; 15:s7=12;
          endcase
        endcase
    end endfunction

    function [3:0] s8; input [5:0] b; integer r,c; begin
        r={b[5],b[0]}; c=b[4:1];
        case(r)
          0: case(c)
            0:s8=13;1:s8=2; 2:s8=8; 3:s8=4; 4:s8=6; 5:s8=15;6:s8=11;7:s8=1;
            8:s8=10;9:s8=9;10:s8=3; 11:s8=14;12:s8=5; 13:s8=0; 14:s8=12;15:s8=7;
          endcase
          1: case(c)
            0:s8=1; 1:s8=15;2:s8=13;3:s8=8; 4:s8=10;5:s8=3; 6:s8=7; 7:s8=4;
            8:s8=12;9:s8=5;10:s8=6; 11:s8=11;12:s8=0; 13:s8=14;14:s8=9; 15:s8=2;
          endcase
          2: case(c)
            0:s8=7; 1:s8=11;2:s8=4; 3:s8=1; 4:s8=9; 5:s8=12;6:s8=14;7:s8=2;
            8:s8=0; 9:s8=6;10:s8=10;11:s8=13;12:s8=15;13:s8=3;14:s8=5; 15:s8=8;
          endcase
          default: case(c)
            0:s8=2; 1:s8=1; 2:s8=14;3:s8=7; 4:s8=4; 5:s8=10;6:s8=8; 7:s8=13;
            8:s8=15;9:s8=12;10:s8=9; 11:s8=0; 12:s8=3; 13:s8=5; 14:s8=6; 15:s8=11;
          endcase
        endcase
    end endfunction

    wire [5:0] b1=in48[47:42], b2=in48[41:36], b3=in48[35:30], b4=in48[29:24];
    wire [5:0] b5=in48[23:18], b6=in48[17:12], b7=in48[11:6],  b8=in48[5:0];

    assign out32 = { s1(b1), s2(b2), s3(b3), s4(b4), s5(b5), s6(b6), s7(b7), s8(b8) };
endmodule

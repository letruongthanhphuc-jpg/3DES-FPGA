// ============================================================================
// 3DES DECRYPT: D(k2) -> E(k1) -> D(k0)
// Input : data_in  (ciphertext)
// Output: data_out (plaintext)
// ============================================================================
module des3_decrypt (
    input         clock,
    input         rst,
    input         select,        // pulse 1 clock để bắt đầu 1 lần 3DES
    input  [63:0] key0,
    input  [63:0] key1,
    input  [63:0] key2,
    input  [63:0] data_in,       // Ciphertext
    output reg [63:0] data_out,  // Plaintext
    output reg        done
);

    // ========================================================================
    //  Key registers
    // ========================================================================
    reg [63:0] k0, k1, k2;

    always @(posedge clock or posedge rst) begin
        if (rst) begin
            k0 <= 64'd0;
            k1 <= 64'd0;
            k2 <= 64'd0;
        end else begin
            k0 <= key0;
            k1 <= key1;
            k2 <= key2;
        end
    end

    // ========================================================================
    //  Wires giữa các stage
    // ========================================================================
    wire [63:0] block0_out;   // output stage 1
    wire [63:0] block1_out;   // output stage 2
    wire [63:0] block2_out;   // output stage 3 (final)

    wire [2:0]  sub_done;     // done từng stage

    // ========================================================================
    //  FSM điều khiển 3 stage
    // ========================================================================
    localparam S_IDLE  = 3'd0,
               S_RUN0  = 3'd1,
               S_WAIT0 = 3'd2,
               S_RUN1  = 3'd3,
               S_WAIT1 = 3'd4,
               S_RUN2  = 3'd5,
               S_WAIT2 = 3'd6;

    reg [2:0] state, nstate;

    // start cho từng block con (nối vào .select)
    reg start0, start1, start2;

    // -------------------------
    //  Next-state & start logic
    // -------------------------
    always @* begin
        // default
        nstate = state;
        start0 = 1'b0;
        start1 = 1'b0;
        start2 = 1'b0;

        case (state)
            // Chờ lệnh start từ trên
            S_IDLE: begin
                if (select) begin
                    nstate = S_RUN0;
                    start0 = 1'b1;           // chạy stage 1
                end
            end

            // Stage 1 đang chạy
            S_RUN0: begin
                if (sub_done[0])            // stage 1 xong
                    nstate = S_WAIT0;
            end

            // 1 clock chờ sau stage 1, rồi kích stage 2
            S_WAIT0: begin
                start1 = 1'b1;              // chạy stage 2
                nstate = S_RUN1;
            end

            // Stage 2 đang chạy
            S_RUN1: begin
                if (sub_done[1])            // stage 2 xong
                    nstate = S_WAIT1;
            end

            // 1 clock chờ sau stage 2, rồi kích stage 3
            S_WAIT1: begin
                start2 = 1'b1;              // chạy stage 3
                nstate = S_RUN2;
            end

            // Stage 3 đang chạy
            S_RUN2: begin
                if (sub_done[2])            // stage 3 xong
                    nstate = S_WAIT2;
            end

            // Chốt kết quả, cho phép vòng mới nếu select=1
            S_WAIT2: begin
                if (select) begin
                    nstate = S_RUN0;
                    start0 = 1'b1;
                end else begin
                    nstate = S_IDLE;
                end
            end

            default: begin
                nstate = S_IDLE;
            end
        endcase
    end

    // -------------------------
    //  State register + output
    // -------------------------
    always @(posedge clock or posedge rst) begin
        if (rst) begin
            state    <= S_IDLE;
            data_out <= 64'd0;
            done     <= 1'b0;
        end else begin
            state <= nstate;

            // done chỉ high 1 clock tại S_WAIT2
            done <= (state == S_WAIT2);

            // chốt ciphertext giải mã xong ở S_WAIT2
            if (state == S_WAIT2)
                data_out <= block2_out;
        end
    end

    // ========================================================================
    //  3 BLOCK DES CON
    //  Encrypt: E(k0) -> D(k1) -> E(k2)
    //  Decrypt: D(k2) -> E(k1) -> D(k0)
    // ========================================================================

    // Stage 1: Decrypt với key2, input là ciphertext
    des_decrypt stage1 (
        .clk          (clock),
        .rst          (rst),
        .select       (start0),
        .ciphertext   (data_in),
        .key          (k2),
        .plaintext_out(block0_out),
        .done         (sub_done[0])
    );

    // Stage 2: Encrypt với key1
    des_encrypt stage2 (
        .clk       (clock),
        .rst       (rst),
        .select    (start1),
        .plaintext (block0_out),
        .key       (k1),
        .dectext   (block1_out),
        .done      (sub_done[1])
    );

    // Stage 3: Decrypt với key0, ra plaintext gốc
    des_decrypt stage3 (
        .clk          (clock),
        .rst          (rst),
        .select       (start2),
        .ciphertext   (block1_out),
        .key          (k0),
        .plaintext_out(block2_out),
        .done         (sub_done[2])
    );

endmodule
